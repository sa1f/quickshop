// pwm_pll.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module pwm_pll (
		input  wire  clk_in_clk,   //   clk_in.clk
		output wire  pwm_clk0_clk, // pwm_clk0.clk
		output wire  pwm_clk1_clk, // pwm_clk1.clk
		output wire  pwm_clk2_clk, // pwm_clk2.clk
		input  wire  rst_in_reset  //   rst_in.reset
	);

	pwm_pll_pll_0 pll_0 (
		.refclk   (clk_in_clk),   //  refclk.clk
		.rst      (rst_in_reset), //   reset.reset
		.outclk_0 (pwm_clk0_clk), // outclk0.clk
		.outclk_1 (pwm_clk1_clk), // outclk1.clk
		.outclk_2 (pwm_clk2_clk), // outclk2.clk
		.locked   ()              // (terminated)
	);

endmodule
