
module pwm_pll (
	clk_in_clk,
	reset_in_reset,
	pwm_clk0_clk,
	pwm_clk1_clk,
	pwm_clk2_clk);	

	input		clk_in_clk;
	input		reset_in_reset;
	output		pwm_clk0_clk;
	output		pwm_clk1_clk;
	output		pwm_clk2_clk;
endmodule
